/*
 * LT24 Test Bench
 * ------------------------
 * By: Thomas Carpenter
 * For: University of Leeds
 * Date: 29th December 2017
 *
 * Description
 * -----------
 * This is a simple test bench module to allow simulation of
 * the LT24 display.
 *
 */

// Timescale indicates unit of delays.
//  `timescale  unit / precision
// Where delays are given as:
//   #unit.precision
//
// For the clock generator in this test bench to work, we must
// stick with a "unit" of 1ns. You may choose the "precision".
//
// e.g for `timescale 1ns/100ps then:
//   #1 = 1ns
//   #1.5 = 1.5ns
//   #1.25 = 1.3ns (rounded to nearest precision)
`timescale 1 ns/100 ps

// Test bench module declaration
//  Always end test bench module names with _tb for clarity
//  There is no port list for a test bench
module LT24Top_tb;

//
// Parameter Declarations
//
localparam NUM_CYCLES = 1000000000;   //Run simulation for NUM_CYCLES clock cycles. (Max 1 billion)
localparam CLOCK_FREQ = 50000000; //Clock frequency

//
// Test Bench Generated Signals
//
reg  clock;
reg  enableLCD;
reg reset;
reg [3:0] valueHr1, valueHr0, valueMin1, valueMin0;
//
// DUT Output Signals
//
wire resetApp;
// LT24 Display Interface
wire        LT24Wr_n;
wire        LT24Rd_n;
wire        LT24CS_n;
wire        LT24RS;
wire        LT24Reset_n;
wire [15:0] LT24Data;
wire        LT24LCDOn;

//
// Device Under Test
//
LT24Top  LT24Top_dut (
   .clock       ( clock ),
   .enableLCD ( reset ),
   .valueHr1(valueHr1),
   .valueHr0(valueHr0),
   .valueMin1(valueMin1),
   .valueMin0(valueMin0),
   .resetApp    ( resetApp    ),   
   .LT24Wr_n    ( LT24Wr_n    ),
   .LT24Rd_n    ( LT24Rd_n    ),
   .LT24CS_n    ( LT24CS_n    ),
   .LT24RS      ( LT24RS      ),
   .LT24Reset_n ( LT24Reset_n ),
   .LT24Data    ( LT24Data    ),
   .LT24LCDOn   ( LT24LCDOn   )
);

initial begin
    $display("%d ns\tSimulation Started",$time);       //Print to console that the simulation has started
    reset = 1'b0;                                      //Start in reset.
    repeat(2) @(posedge clock);                        //Wait for a couple of clock cycles
    reset = 1'b1;                                      //Then clear the reset signal.
    wait(resetApp === 1'b0);                           //Wait until the resetApp signal is zero.
    $display("%d ns\tInitialisation Successful",$time);  //Print to console that initialisation of the display is complete.
	$display("Initialisation verified. LCD ready to take values"); 				// Initialisation verified.
	//once complete assign time values
	valueHr1 = 4'd0;
	valueHr0 = 4'd9;
	valueMin1 = 4'd0;
	valueMin0 = 4'd15;
	
end


//
//Clock generator + simulation time limit.
//

initial begin
    clock = 1'b0; //Initialise the clock to zero.
end

//Next we convert our clock period to nanoseconds and half it
//to work out how long we must delay for each half clock cycle
real HALF_CLOCK_PERIOD = (1000000000.0 / $itor(CLOCK_FREQ)) / 2.0;

//Now generate the clock
integer half_cycles = 0;
always begin
    //Generate the next half cycle of clock
    #(HALF_CLOCK_PERIOD);          //Delay for half a clock period.
    clock = ~clock;                //Toggle the clock
    half_cycles = half_cycles + 1; //Increment the counter
    //$monitor("NUM_CYCLES=%d",half_cycles);
    //Check if enough half clock cycle
    if (half_cycles == (2*NUM_CYCLES)) begin 
        //Once the number of cycles has been reached
		half_cycles = 0; 		   //Reset half cycles, so if we resume running with "run -all", we perform another chunk.
		$monitor("NUM_CYCLES=%d",NUM_CYCLES);
		$display("%d ns\tInitialisation in progress",$time);
        $stop;                     //Break the simulation
		
        //Note: We can continue the simulation after this breakpoint using "run -continue" or "run x ns" or "run -all" in modelsim.
    end
end
endmodule
